library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity LCDDriver is
  generic (
    
  );
  port (
  );
end entity;

architecture rtl of LCDDriver is
begin
end architecture;