library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;

entity DisplayDriverALU4_4FP is
    port (
        i_CLK       : in  std_logic;
        i_Number    : in  std_logic_vector(7 downto 0);
        o_Displays  : out std_logic_vector(3 downto 0);
        o_Segments  : out std_logic_vector(6 downto 0);
        o_DispPoint : out std_logic
    );
end entity DisplayDriverALU4_4FP;

architecture rtl of DisplayDriverALU4_4FP is
    
    component BCDTo7Segs is
        port (
            i_DispPoint       : in  std_logic;                     --Display point enable
            i_ChipEn          : in  std_logic;                     --Chip enable (works with PNP transistors)
            i_Number          : in  std_logic_vector(3 downto 0);  --Number that will be displayed
            o_DisplaySegments : out std_logic_vector(6 downto 0);  --Display segments vector
            o_DispEnable      : out std_logic;                     --Out pin to enable the display (works with i_ChipEn)
            o_DispPoint       : out std_logic                      --Turns up or down the display point (works with i_DispPoint)
        );
    end component BCDTo7Segs;
    
    constant DISP_NEGATIVE_SIGN       : std_logic_vector(6 downto 0) := "0111111";
    constant DISP_POSITIVE_SIGN       : std_logic_vector(6 downto 0) := "1111111";
	signal r_Sel   					  : std_logic_vector(1 downto 0) := "00";
	signal r_Show  					  : std_logic_vector(3 downto 0) := "0000";
    signal r_IntPNumber, r_DecPNumber : std_logic_vector(3 downto 0);
    signal r_Segs1, r_Segs2           : std_logic_vector(6 downto 0);
    signal r_SegsConn1, r_SegsConn2   : std_logic_vector(6 downto 0);
    signal r_NumberSign               : std_logic;
	signal r_Count					  : integer range 0 to 100000;

begin
    
    DisplayDecoder1 : BCDTo7Segs port map (
        i_DispPoint       => '1',
        i_ChipEN          => '1',
        i_Number          => r_IntPNumber,
        o_DisplaySegments => r_SegsConn1,
        o_DispPoint       => o_DispPoint
    );

    DisplayDecoder2 : BCDTo7Segs port map (
        i_DispPoint        => '0',
        i_ChipEN           => '1',
        i_Number           => r_DecPNumber,
        o_DisplaySegments   => r_SegsConn2
    );

    clkCount : process(i_CLK)
    begin
        if rising_edge(i_CLK) then
            if r_Count < 10 then --100000
                r_Count <= r_Count + 1;
            else 
                r_Sel <= r_Sel + 1;
                r_Count <= 0;
            end if;
        end if;
    end process;

    ShowDisplays : process(r_Sel, r_NumberSign, r_SegsConn1, r_SegsConn2, r_Segs1, r_Segs2, r_Show)
    begin
        r_Segs1 <= r_SegsConn1;
        r_Segs2 <= r_SegsConn2;
        case r_Sel is
            when "00" => 
                r_Show <= "1110";
            when "01" =>
                r_Show <= "1101";
            when "10" =>
                r_Show <= "1011";
            when "11" =>
                r_Show <= "0111";
            when others =>
                r_Show <= "1111";
        end case;
        
        if r_NumberSign = '1' then
            r_Segs1 <= r_Segs1 + 1;
            r_Segs1 <= not r_Segs1; 
            r_Segs2 <= r_Segs2 + 1;
            r_Segs2 <= not r_Segs2; 
        end if;

        case r_Show is
            when "1101" => --3
                o_Segments <= r_Segs2;
            when "1011" => --2
                o_Segments <= r_Segs1;
            when "0111" => --1
                case r_NumberSign is
                    when '1' =>
                        o_Segments <= DISP_NEGATIVE_SIGN;
                    when others =>
                        o_Segments <= DISP_POSITIVE_SIGN;
                end case;
            when others =>
                o_Segments <= "1111111";
        end case;    
    end process;
    
    r_IntPNumber <= i_Number(7 downto 4);

    r_DecPNumber <= i_Number(3 downto 0);

    o_Displays <= r_Show;

    r_NumberSign <= i_Number(7);
    
end architecture rtl;